`ifndef FULL_FUNCTION_ARITHMETIC_LOGICAL_UNIT_32BIT_V
`define FULL_FUNCTION_ARITHMETIC_LOGICAL_UNIT_32BIT_V

module ALU32 (
    input  wire [ 3:0] ctl,
    input  wire [31:0] rs1,
    input  wire [31:0] rs2,
    output wire [31:0] rd,
);

endmodule

`endif 