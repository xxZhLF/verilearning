`ifndef ADD_32BIT_FLOAT_V
`define ADD_32BIT_FLOAT_V

module Add32F(
    input  wire [31:0] op1,
    input  wire [31:0] op2,
    output wire [31:0] sum
);



endmodule

`endif 