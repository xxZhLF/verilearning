`ifndef MICROARCHITECTURE_SINGLE_CYCLE_V
`define MICROARCHITECTURE_SINGLE_CYCLE_V

module MicroarchSC (
    input wire rst;
    input wire clk;
);
    
endmodule

`endif 