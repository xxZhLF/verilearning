`include "Add64.v"
`include "Shift.v"

module MulBT32S(
    input  wire [31:0] op1,
    input  wire [31:0] op2,
    output wire [63:0] res
);

endmodule

module BoothEncoding (
    input  wire[ 2:0] grp,  // Group of 3-bit 
    input  wire[ 2:0] gid,  // Index of Group
    input  wire[31:0] op1,  // Multiplier
    output wire[63:0] pp    // Partial Product
);

    wire       sb;
    wire [8:0] nb;

    assign {sb, nb} = ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd0}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd1}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd2}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd3}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd4}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd5}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd6}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b000} | ~|{grp ^ 3'b111}) & ~|{gid ^ 3'd7}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd0}) ? {1'b0, 8'h00} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd1}) ? {1'b0, 8'h02} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd2}) ? {1'b0, 8'h04} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd3}) ? {1'b0, 8'h06} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd4}) ? {1'b0, 8'h08} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd5}) ? {1'b0, 8'h0A} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd6}) ? {1'b0, 8'h0C} : 
                      ((~|{grp ^ 3'b001} | ~|{grp ^ 3'b010}) & ~|{gid ^ 3'd7}) ? {1'b0, 8'h0E} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd0}) ? {1'b0, 8'h02} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd1}) ? {1'b0, 8'h04} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd2}) ? {1'b0, 8'h06} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd3}) ? {1'b0, 8'h08} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd4}) ? {1'b0, 8'h0A} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd5}) ? {1'b0, 8'h0C} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd6}) ? {1'b0, 8'h0E} : 
                      ((~|{grp ^ 3'b011}                   ) & ~|{gid ^ 3'd7}) ? {1'b0, 8'h10} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd0}) ? {1'b1, 8'h02} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd1}) ? {1'b1, 8'h04} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd2}) ? {1'b1, 8'h06} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd3}) ? {1'b1, 8'h08} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd4}) ? {1'b1, 8'h0A} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd5}) ? {1'b1, 8'h0C} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd6}) ? {1'b1, 8'h0E} : 
                      ((~|{grp ^ 3'b100}                   ) & ~|{gid ^ 3'd7}) ? {1'b1, 8'h10} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd0}) ? {1'b1, 8'h00} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd1}) ? {1'b1, 8'h02} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd2}) ? {1'b1, 8'h04} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd3}) ? {1'b1, 8'h06} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd4}) ? {1'b1, 8'h08} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd5}) ? {1'b1, 8'h0A} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd6}) ? {1'b1, 8'h0C} : 
                      ((~|{grp ^ 3'b101} | ~|{grp ^ 3'b110}) & ~|{gid ^ 3'd7}) ? {1'b1, 8'h0E} : {1'bZ, 8'hZZ};

    ShiftL64 shift(
        .n(nb),
        .in({32'h0, op1}),
        .out(pp)
    );

    // 根据符号判断：是将原码转换为补码，还是将补码转换为原码
    
endmodule