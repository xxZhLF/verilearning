`timescale 1ps/1ps 

module MicroarchSC_tb(
    // None
);

endmodule