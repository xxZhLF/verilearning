`include "AdderHF1bit.v"

module AdderHF1bit_tb (
    // None
);
    initial begin
        $display("Hello World!");
        $finish;
    end
    
    // AdderHF1bit adder();

endmodule