`ifndef MICROARCHITECTURE_SINGLE_CYCLE_V
`define MICROARCHITECTURE_SINGLE_CYCLE_V

`include "../IPs_shared/universal4inc.v"
`include "../0x0101_ALU32FF/CtlALU.v"
`include "../0x0200_REGs3P/RegName.v"
`include "../0x0300_PC/PCIM.v"
`include "../0x0400_Decoder/RV32I.v"
`include "../0x0400_Decoder/RV32M.v"
`include "../0x0500_Mem/MemIO.v"

`define DATA_ST `MM_ENB_W
`define DATA_LD `MM_ENB_R

module MicroarchiSC (
    input  wire        rst,
    input  wire        clk_LF,
    input  wire        clk_HF,
    input  wire [31:0] instr,
    input  wire [31:0] dataI,
    output wire [31:0] dataO,
    output wire        store_or_load,
    output wire [ 1:0] width_of_data,
    output wire [31:0] locat_of_data,
    output wire [31:0] where_is_instr
);

    reg clk_UC; /* UnConventional */
    always @(posedge clk_LF) 
        clk_UC <= rst ? 1'b1 : ~clk_UC;

    wire [ 1:0] pc_mode;
    wire [31:0] pc_offset;
    wire [31:0] pc_target;
    wire [31:0] pc_addr;
    wire [31:0] pc_addr_nxt;
    PC pc(
        .rst(rst),
        .clk(clk_UC),
        .mode(pc_mode),
        .offset(pc_offset),
        .target(pc_target),
        .addr(pc_addr),
        .addr_ret(pc_addr_nxt)
    );

    wire        rf_en4w;
    wire [ 4:0] rf_wA;
    wire [31:0] rf_wD;
    wire [ 4:0] rf_r0A, rf_r1A;
    wire [31:0] rf_r0D, rf_r1D;
    REGs3P rf(
        .clk(clk_HF),
        .en4w(rf_en4w),
        .addr_w(rf_wA),
        .data_i(rf_wD),
        .addr_r0(rf_r0A),
        .data_o0(rf_r0D),
        .addr_r1(rf_r1A),
        .data_o1(rf_r1D)
    );

    wire [15:0] alu_ctl;
    wire [31:0] alu_op1;
    wire [31:0] alu_op2;
    wire [31:0] alu_res;
    ALU32FF alu(
        .ctl(alu_ctl),
        .op1(alu_op1),
        .op2(alu_op2),
        .res(alu_res)
    );

    wire [31:0] decoder_instr;
    wire [ 6:0] decoder_op;
    wire [ 4:0] decoder_rs1;
    wire [ 4:0] decoder_rs2;
    wire [ 4:0] decoder_rd;
    wire [ 9:0] decoder_func;
    wire [31:0] decoder_imm;
    Decoder decoder(
        .instr(decoder_instr),
        .op(decoder_op),
        .rs1(decoder_rs1),
        .rs2(decoder_rs2),
        .rd(decoder_rd),
        .func(decoder_func),
        .imm(decoder_imm)
    );

    wire [31:0] c2t_1C, c2t_2C;
    wire [31:0] c2t_1T, c2t_2T;
    CTC32 c2t_1(
        .C(c2t_1C),
        .T(c2t_1T)
    ), c2t_2(
        .C(c2t_2C),
        .T(c2t_2T)
    );

    wire [31:0] c2t_IC;
    wire [31:0] c2t_IT;
    CTC32 c2t_I(
        .C(c2t_IC),
        .T(c2t_IT)
    );

    wire [31:0] t2c_T;
    wire [31:0] t2c_C;
    TCC32 t2c(
        .T(t2c_T),
        .C(t2c_C)
    );

    parameter HB = 32 +  1 +  2 + 32 +  1 
                 +  5 + 32 +  5 +  5 +  2 
                 + 32 + 32 + 16 + 32 + 32 
                 + 32 + 32 + 32 + 32 ;
    wire [HB-1 : 0] I2Hub, Hub2O;
    assign {
    /* No.18: 32-Bit */ dataO, /*         [388:357] Date Wrote to Memory                         */
    /* No.17:  1-Bit */ store_or_load, /* [    356] Signal of Memory Read/Write                  */
    /* No.16:  2-Bit */ width_of_data, /* [355:354] Size of Date in Memory to Read/Write         */
    /* No.15: 32-Bit */ locat_of_data, /* [353:322] Address of Memory to Read/Write              */
    /* No.14:  1-Bit */ rf_en4w, /*       [    321] Write Signal of Destination Register         */
    /* No.13:  5-Bit */ rf_wA, /*         [320:316] Address of Destination Register              */
    /* No.12: 32-Bit */ rf_wD, /*         [315:284] Value Write to Destination Register          */
    /* No.11:  5-Bit */ rf_r0A, /*        [283:279] Address of Source Register 1                 */
    /* No.10:  5-Bit */ rf_r1A, /*        [278:274] Address of Source Register 2                 */
    /* No.9:   2-Bit */ pc_mode, /*       [273:272] Mode of PC                                   */
    /* No.8:  32-Bit */ pc_offset, /*     [271:240] Offset Add to PC                             */
    /* No.7:  32-Bit */ pc_target, /*     [239:208] Target Write to PC                           */
    /* No.6:  16-Bit */ alu_ctl, /*       [207:192] Control Signal of ALU                        */
    /* No.5:  32-Bit */ alu_op1, /*       [191:160] OP1 of ALU                                   */
    /* No.4:  32-Bit */ alu_op2, /*       [159:128] OP2 of ALU                                   */
    /* No.3:  32-Bit */ c2t_1C, /*        [127: 96] 2'complement (Converted to True Code as OP1) */
    /* No.2:  32-Bit */ c2t_2C, /*        [ 95: 64] 2'complement (Converted to True Code as OP2) */
    /* No.1:  32-Bit */ c2t_IC, /*        [ 63: 32] 2'complement (Converted to True Code as IMM) */
    /* No.0:  32-Bit */ t2c_T /*          [ 31:  0] RES of True Code (Converted to 2'complement) */                /* No.18: 32-Bit  */ /* No.17: 1-Bit  */ /* No.16: 2-Bit  */ /* No.15: 32-Bit  */ /* No.14: 1-Bit */ /* No.13: 5-Bit  */ /* No.12: 32-Bit                     */ /* No.11: 5-Bit   */ /* No.10: 5-Bit   */ /* No.9: 2-Bit */ /* No.8: 32-Bit                                   */ /* No.7: 32-Bit  */ /* No.6: 16-Bit     */ /* No.5: 32-Bit            */ /* No.4: 32-Bit                  */ /* No.3: 32-Bit        */ /* No.2: 32-Bit        */ /* No.1: 32-Bit        */ /* No.0: 32-Bit                               */
    } = Hub2O; assign I2Hub = `isEQ(decoder_op, `INSTR_TYP_R)     ? `isEQ(decoder_func, `R_TYP_FC_ADD)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_SUB)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SUB,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_SLL)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLL,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_SRL)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SRL,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_SRA)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SRA,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_SLT)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLT,  /* | */ c2t_1T,               /* | */ c2t_2T,                     /* | */ rf_r0D,           /* | */ rf_r1D,           /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_SLTU)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLTU, /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_AND)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_AND,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_OR)       ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_OR,   /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_XOR)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_XOR,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_MUL)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_MUL,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_MULH)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_MUL,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_MULHU)    ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_MUL,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_MULHSU )  ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_MUL,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_DIV)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ t2c_C,                          /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_DIV,  /* | */ {1'b0, c2t_1T[30:0]}, /* | */ {1'b0, c2t_2T[30:0]},       /* | */ rf_r0D,           /* | */ rf_r1D,           /* | */ {32{1'bZ}},       /* | */ {rf_r0D[31] ^ rf_r1D[31], alu_res[30:0]} /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_REM)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_REM,  /* | */ {1'b0, c2t_1T[30:0]}, /* | */ {1'b0, c2t_2T[30:0]},       /* | */ rf_r0D,           /* | */ rf_r1D,           /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_DIVU)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_DIV,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `R_TYP_FC_REMU)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_REM,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_I)     ? `isEQ(decoder_func, `I_TYP_FC_ADDI)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_SLTI)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLT,  /* | */ c2t_1T,               /* | */ c2t_IT,                     /* | */ rf_r0D,           /* | */ {32{1'bZ}},       /* | */ decoder_imm,      /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_SLTIU)    ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLTU, /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_ANDI)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_AND,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_ORI)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_OR,   /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_XORI)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_XOR,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_SLLI)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLL,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_SRLI)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SRL,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I_TYP_FC_SRAI)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SRA,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_S)     ? `isEQ(decoder_func, `S_TYP_FC_SB)       ? {/* | */ rf_r1D,      /* | */ `DATA_ST,   /* | */ `MW_Byte,   /* | */ alu_res,     /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `S_TYP_FC_SH)       ? {/* | */ rf_r1D,      /* | */ `DATA_ST,   /* | */ `MW_Half,   /* | */ alu_res,     /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `S_TYP_FC_SW)       ? {/* | */ rf_r1D,      /* | */ `DATA_ST,   /* | */ `MW_Word,   /* | */ alu_res,     /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_B)     ? `isEQ(decoder_func, `B_TYP_FC_BEQ)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ {5{1'bZ}},   /* | */ {5{1'bZ}},   /* | */ `BRANCH,  /* | */ `isEQ(rf_r0D, rf_r1D) ? decoder_imm : 32'd4, /* | */ {32{1'bZ}}, /* | */ {16{1'bZ}},    /* | */ {32{1'bZ}},           /* | */ {32{1'bZ}},                 /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `B_TYP_FC_BEN)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ {5{1'bZ}},   /* | */ {5{1'bZ}},   /* | */ `BRANCH,  /* | */ `isEQ(rf_r0D, rf_r1D) ? 32'd4 : decoder_imm, /* | */ {32{1'bZ}}, /* | */ {16{1'bZ}},    /* | */ {32{1'bZ}},           /* | */ {32{1'bZ}},                 /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `B_TYP_FC_BLT)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `BRANCH,  /* | */            alu_res[0] ? decoder_imm : 32'd4, /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLT,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `B_TYP_FC_BGE)      ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `BRANCH,  /* | */            alu_res[0] ? 32'd4 : decoder_imm, /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLT,  /* | */ rf_r0D,               /* | */ rf_r1D,                     /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `B_TYP_FC_BLTU)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `BRANCH,  /* | */            alu_res[0] ? decoder_imm : 32'd4, /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLTU, /* | */ c2t_1T,               /* | */ c2t_2T,                     /* | */ rf_r0D,           /* | */ rf_r1D,           /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `B_TYP_FC_BGEU)     ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'bZ,      /* | */ {5{1'bZ}},  /* | */ {32{1'bZ}},                     /* | */ decoder_rs1, /* | */ decoder_rs2, /* | */ `BRANCH,  /* | */            alu_res[0] ? 32'd4 : decoder_imm, /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_SLTU, /* | */ c2t_1T,               /* | */ c2t_2T,                     /* | */ rf_r0D,           /* | */ rf_r1D,           /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* ========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_U)     ?                                    1'b1 ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ decoder_imm,                    /* | */ {5{1'bZ}},   /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ {16{1'bZ}},    /* | */ {32{1'bZ}},           /* | */ {32{1'bZ}},                 /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_J)     ?                                    1'b1 ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ pc_addr_nxt,                    /* | */ {5{1'bZ}},   /* | */ {5{1'bZ}},   /* | */ `UCJUMP,  /* | */ {32{1'bZ}},                                  /* | */ alu_res,    /* | */ `ALU_CTL_ADD,  /* | */ pc_addr,              /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_I12LD) ? `isEQ(decoder_func, `I12LD_TYP_FC_LB)   ? {/* | */ {32{1'bZ}},  /* | */ `DATA_LD,   /* | */ `MW_Byte,   /* | */ alu_res,     /* | */ 1'b1,      /* | */ decoder_rd, /* | */ {{24{dataI[ 7]}}, dataI[ 7:0]}, /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I12LD_TYP_FC_LH)   ? {/* | */ {32{1'bZ}},  /* | */ `DATA_LD,   /* | */ `MW_Half,   /* | */ alu_res,     /* | */ 1'b1,      /* | */ decoder_rd, /* | */ {{16{dataI[15]}}, dataI[15:0]}, /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I12LD_TYP_FC_LW)   ? {/* | */ {32{1'bZ}},  /* | */ `DATA_LD,   /* | */ `MW_Word,   /* | */ alu_res,     /* | */ 1'b1,      /* | */ decoder_rd, /* | */ dataI,                          /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I12LD_TYP_FC_LBU)  ? {/* | */ {32{1'bZ}},  /* | */ `DATA_LD,   /* | */ `MW_Byte,   /* | */ alu_res,     /* | */ 1'b1,      /* | */ decoder_rd, /* | */ {24'b0, dataI[ 7:0]},           /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : 
                                                                    `isEQ(decoder_func, `I12LD_TYP_FC_LBU)  ? {/* | */ {32{1'bZ}},  /* | */ `DATA_LD,   /* | */ `MW_Byte,   /* | */ alu_res,     /* | */ 1'b1,      /* | */ decoder_rd, /* | */ {16'b0, dataI[15:0]} ,          /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_I12JR) ? `isEQ(decoder_func, `I12JR_TYP_FC_JALR) ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ pc_addr_nxt,                    /* | */ decoder_rs1, /* | */ {5{1'bZ}},   /* | */ `UCJUMP,  /* | */ {32{1'bZ}},                                  /* | */ alu_res,    /* | */ `ALU_CTL_ADD,  /* | */ rf_r0D,               /* | */ decoder_imm,                /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} :
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */
                              `isEQ(decoder_op, `INSTR_TYP_I20PC) ?                                    1'b1 ? {/* | */ {32{1'bZ}},  /* | */ 1'bZ,       /* | */ 2'bZZ,      /* | */ {32{1'bZ}},  /* | */ 1'b1,      /* | */ decoder_rd, /* | */ alu_res,                        /* | */ {5{1'bZ}},   /* | */ {5{1'bZ}},   /* | */ `NORMAL,  /* | */ {32{1'bZ}},                                  /* | */ {32{1'bZ}}, /* | */ `ALU_CTL_ADD,  /* | */ pc_addr,              /* | */ {decoder_imm[19:0], 12'b0}, /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}},       /* | */ {32{1'bZ}}                               /* | */} : {HB{1'bZ}} : {HB{1'bZ}};
                                                                  /* =========================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================================== */


    assign decoder_instr = instr;
    assign where_is_instr = rst ? 32'h800 : pc_addr;

    reg [HB-1 : 0] __Hub__;
    assign Hub2O = __Hub__;
    always @(negedge rst or posedge clk_LF) begin
        if (rst) begin 
            __Hub__[273:272] <= `UCJUMP; /* PC Mode   */
            __Hub__[239:208] <= 32'h800; /* PC Target */
        end else begin 
            __Hub__ <= I2Hub;
        end
    end

`define DBG_TRACE_LOG_ENABLE
`ifndef DBG_TRACE_LOG_ENABLE
`else

    reg [31:0] cnt;
    always @(posedge clk_UC) 
        cnt <= rst ? 0'b0 : cnt + 32'b1;

    reg [ 6:0] DBG_decoder_op;
    reg [ 9:0] DBG_decoder_func;
    reg [31:0] DBG_decoder_imm;

    always @(posedge clk_LF) begin
        if (rst) begin
        end else begin
            DBG_decoder_op   <= decoder_op;
            DBG_decoder_func <= decoder_func;
            DBG_decoder_imm  <= decoder_imm;
            if (clk_UC) begin
            end else begin
                DBG_detail_of_instr_exec(cnt,
                                         pc_addr,
                                         decoder_instr, 
                                         DBG_decoder_op,   /* As output of module, transit by debug register */
                                         DBG_decoder_func, /* As output of module, transit by debug register */
                                         DBG_decoder_imm,  /* As output of module, transit by debug register */
                                         rf_r0A, rf_r0D,   /* As  input of module, transit by Hub */
                                         rf_r1A, rf_r1D,   /* As  input of module, transit by Hub */
                                         rf_wA,  rf_wD);   /* As  input of module, transit by Hub */
            end
        end
    end

    task DBG_detail_of_instr_exec(
        input [31:0] idx,
        input [31:0] pc,
        input [31:0] instr,
        input [ 6:0] op,
        input [ 9:0] func,
        input [31:0] imm,
        input [ 4:0] rs1_addr,
        input [31:0] rs1_data,
        input [ 4:0] rs2_addr, 
        input [31:0] rs2_data,
        input [ 4:0]  rd_addr,
        input [31:0]  rd_data
    ); begin
        case (op)
            `INSTR_TYP_R: begin
                case (func)
                    `R_TYP_FC_ADD:      $display("No.%03d ADD:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_SUB:      $display("No.%03d SUB:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_SLL:      $display("No.%03d SLL:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_SLT:      $display("No.%03d SLT:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_SLTU:     $display("No.%03d SLTU:   @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_XOR:      $display("No.%03d XOR:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_SRL:      $display("No.%03d SRL:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_SRA:      $display("No.%03d SRA:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_OR:       $display("No.%03d OR:     @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_AND:      $display("No.%03d AND:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_MUL:      $display("No.%03d MUL:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_MULH:     $display("No.%03d MULH:   @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_MULHSU:   $display("No.%03d MULHSU: @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_MULHU:    $display("No.%03d MULHU:  @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_DIV:      $display("No.%03d DIV:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_DIVU:     $display("No.%03d DIVU:   @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_REM:      $display("No.%03d REM:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    `R_TYP_FC_REMU:     $display("No.%03d REMU:   @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, rd  is x%-2d", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, rd_addr);
                    default: $display("*[ERROR]@INSTR_TYP_R Func=%b ", func);
                endcase
            end 
            `INSTR_TYP_I: begin
                case (func)
                    `I_TYP_FC_ADDI:     $display("No.%03d ADDI:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_SLTI:     $display("No.%03d SLTI:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_SLTIU:    $display("No.%03d SLTIU:  @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_XORI:     $display("No.%03d XORI:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_ORI:      $display("No.%03d ORI:    @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_ANDI:     $display("No.%03d ANDI:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_SLLI:     $display("No.%03d SLLI:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_SRLI:     $display("No.%03d SRLI:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I_TYP_FC_SRAI:     $display("No.%03d SRAI:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    default: $display("*[ERROR]@INSTR_TYP_I Func=%b ", func);
                endcase
            end 
            `INSTR_TYP_S: begin
                case (func)
                    `S_TYP_FC_SB:       $display("No.%03d SB:     @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    `S_TYP_FC_SH:       $display("No.%03d SH:     @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    `S_TYP_FC_SW:       $display("No.%03d SW:     @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    default: $display("*[ERROR]@INSTR_TYP_S Func=%b ", func);
                endcase
            end 
            `INSTR_TYP_B: begin
                case (func)
                    `B_TYP_FC_BEQ:      $display("No.%03d BEQ:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    `B_TYP_FC_BEN:      $display("No.%03d BNE:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    `B_TYP_FC_BLT:      $display("No.%03d BLT:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    `B_TYP_FC_BGE:      $display("No.%03d BGE:    @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    `B_TYP_FC_BLTU:     $display("No.%03d BLTU:   @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    `B_TYP_FC_BGEU:     $display("No.%03d BGEU:   @[%08H] rs1 is x%-2d=0x%08H, rs2 is x%-2d=0x%08H, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rs2_addr, rs2_data, imm);
                    default: $display("*[ERROR]@INSTR_TYP_B Func=%b ", func);
                endcase
            end 
            `INSTR_TYP_U: begin
                                        $display("No.%03d LUI:    @[%08H] rd  is x%-2d, imm is 0x%05H", idx, pc, rd_addr, imm);
            end 
            `INSTR_TYP_J: begin
                                        $display("No.%03d JAL:    @[%08H] rd  is x%-2d, imm is 0x%05H", idx, pc, rd_addr, imm);
            end 
            `INSTR_TYP_I12LD: begin
                case (func) 
                    `I12LD_TYP_FC_LB:   $display("No.%03d LB:     @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I12LD_TYP_FC_LH:   $display("No.%03d LH:     @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I12LD_TYP_FC_LW:   $display("No.%03d LW:     @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I12LD_TYP_FC_LBU:  $display("No.%03d LBU:    @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    `I12LD_TYP_FC_LHU:  $display("No.-03d LHU:    @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    default: $display("*[ERROR]@INSTR_TYP_I12LD Func=%b ", func);
                endcase
            end
            `INSTR_TYP_I12JR: begin
                case (func) 
                    `I12JR_TYP_FC_JALR: $display("No.%-3d JALR:   @[%08H] rs1 is x%-2d=0x%08H, rd  is x%-2d, imm is 0x%08H", idx, pc, rs1_addr, rs1_data, rd_addr, imm);
                    default: $display("*[ERROR]@INSTR_TYP_I12JR Func=%b ", func);
                endcase
            end
            `INSTR_TYP_I20PC: begin
                                        $display("No.%-3d AUIPC:  @[%08H] rd  is x%-2d, imm is 0x%05H", idx, pc, rd_addr, imm);
            end
            default: begin
                $display("*[ERROR] Machine Code is instr=%08H, @[%08H]", instr, pc);
            end
        endcase
    end endtask

`endif /* DBG_TRACE_LOG_ENABLE */

endmodule

`endif 