// `define ADD_DEBUG_ON

module AdderLC32bit (
    input  wire [31:0] op1,
    input  wire [31:0] op2,
    input  wire        cin,
    output wire [31:0] sum,
    output wire        cout
`ifdef ADD_DEBUG_ON
  , output wire [31:0] debug
`endif 
);

    // assign {cout, sum} = op1 + op2 + {24'h000000, 7'b00000000, cin};

    wire [31:0] P, G;
    GrpPG grpPG(
        .op1(op1),
        .op2(op2),
        .P(P),
        .G(G)
    );

    wire [31:0] cinner;
    Carry carry(
        .P(P),
        .G(G),
        .cin(cin),
        .cinner(cinner),
        .cout(cout)
    );

    generate
        for (genvar i = 0; i < 32; ++i) begin
            // assign sum[i] = op1[i] ^ op2[i] ^ cinner[i];
            reg useless;
            AdderFL1bit adderFL1bit(
                .op1(op1[i]),
                .op2(op2[i]),
                .cin(cinner[i]),
                .sum(sum[i]),
                .cout(useless)
            );
        end        
    endgenerate

`ifdef ADD_DEBUG_ON
    assign debug = cinner;
    // assign debug = P;
    // assign debug = G;
`endif 

endmodule

module Carry(
    input  wire [31:0] P,
    input  wire [31:0] G,
    input  wire        cin,
    output wire [31:0] cinner,
    output wire        cout
);

    assign {cout, cinner} = {
        /* cout       */ |{ &{G[31]},
                            &{G[30], P[31]},
                            &{G[29], P[30], P[31]},
                            &{G[28], P[29], P[30], P[31]},
                            &{G[27], P[28], P[29], P[30], P[31]},
                            &{G[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]}, 
                            &{G[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]}, 
                            &{G[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], P[31], cin}},
        // /* cout       */ 1'b0,
        /* cinner[31] */ |{ &{G[30]},
                            &{G[29], P[30]},
                            &{G[28], P[29], P[30]},
                            &{G[27], P[28], P[29], P[30]},
                            &{G[26], P[27], P[28], P[29], P[30]},
                            &{G[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]}, 
                            &{G[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]}, 
                            &{G[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], P[30], cin}},
        // /* cinner[31] */ 1'b0,
        /* cinner[30] */ |{ &{G[29]},
                            &{G[28], P[29]},
                            &{G[27], P[28], P[29]},
                            &{G[26], P[27], P[28], P[29]},
                            &{G[25], P[26], P[27], P[28], P[29]},
                            &{G[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]}, 
                            &{G[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]}, 
                            &{G[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], P[29], cin}},
        // /* cinner[30] */ 1'b0,
        /* cinner[29] */ |{ &{G[28]},
                            &{G[27], P[28]},
                            &{G[26], P[27], P[28]},
                            &{G[25], P[26], P[27], P[28]},
                            &{G[24], P[25], P[26], P[27], P[28]},
                            &{G[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[22], P[23], P[24], P[25], P[26], P[27], P[28]}, 
                            &{G[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]}, 
                            &{G[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], P[28], cin}},
        // /* cinner[29] */ 1'b0,
        /* cinner[28] */ |{ &{G[27]},
                            &{G[26], P[27]},
                            &{G[25], P[26], P[27]},
                            &{G[24], P[25], P[26], P[27]},
                            &{G[23], P[24], P[25], P[26], P[27]},
                            &{G[22], P[23], P[24], P[25], P[26], P[27]}, 
                            &{G[21], P[22], P[23], P[24], P[25], P[26], P[27]}, 
                            &{G[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], P[27], cin}},
        // /* cinner[28] */ 1'b0,
        /* cinner[27] */ |{ &{G[26]},
                            &{G[25], P[26]},
                            &{G[24], P[25], P[26]},
                            &{G[23], P[24], P[25], P[26]},
                            &{G[22], P[23], P[24], P[25], P[26]}, 
                            &{G[21], P[22], P[23], P[24], P[25], P[26]}, 
                            &{G[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], P[26], cin}},
        // /* cinner[27] */ 1'b0,
        /* cinner[26] */ |{ &{G[25]},
                            &{G[24], P[25]},
                            &{G[23], P[24], P[25]},
                            &{G[22], P[23], P[24], P[25]}, 
                            &{G[21], P[22], P[23], P[24], P[25]}, 
                            &{G[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], P[25], cin}},
        // /* cinner[26] */ 1'b0,
        /* cinner[25] */ |{ &{G[24]},
                            &{G[23], P[24]},
                            &{G[22], P[23], P[24]}, 
                            &{G[21], P[22], P[23], P[24]}, 
                            &{G[20], P[21], P[22], P[23], P[24]},
                            &{G[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], P[24], cin}},
        // /* cinner[25] */ 1'b0,
        /* cinner[24] */ |{ &{G[23]},
                            &{G[22], P[23]}, 
                            &{G[21], P[22], P[23]}, 
                            &{G[20], P[21], P[22], P[23]},
                            &{G[19], P[20], P[21], P[22], P[23]},
                            &{G[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], P[23], cin}},
        // /* cinner[24] */ 1'b0,
        /* cinner[23] */ |{ &{G[22]}, 
                            &{G[21], P[22]}, 
                            &{G[20], P[21], P[22]},
                            &{G[19], P[20], P[21], P[22]},
                            &{G[18], P[19], P[20], P[21], P[22]},
                            &{G[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], P[22], cin}},
        // /* cinner[23] */ 1'b0,
        /* cinner[22] */ |{ &{G[21]}, 
                            &{G[20], P[21]},
                            &{G[19], P[20], P[21]},
                            &{G[18], P[19], P[20], P[21]},
                            &{G[17], P[18], P[19], P[20], P[21]},
                            &{G[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], P[21], cin}},
        // /* cinner[22] */ 1'b0,
        /* cinner[21] */ |{ &{G[20]},
                            &{G[19], P[20]},
                            &{G[18], P[19], P[20]},
                            &{G[17], P[18], P[19], P[20]},
                            &{G[16], P[17], P[18], P[19], P[20]},
                            &{G[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], P[20], cin}},
        // /* cinner[21] */ 1'b0,
        /* cinner[20] */ |{ &{G[19]},
                            &{G[18], P[19]},
                            &{G[17], P[18], P[19]},
                            &{G[16], P[17], P[18], P[19]},
                            &{G[15], P[16], P[17], P[18], P[19]},
                            &{G[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], P[19], cin}},
        // /* cinner[20] */ 1'b0,
        /* cinner[19] */ |{ &{G[18]},
                            &{G[17], P[18]},
                            &{G[16], P[17], P[18]},
                            &{G[15], P[16], P[17], P[18]},
                            &{G[14], P[15], P[16], P[17], P[18]},
                            &{G[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], P[18], cin}},
        // /* cinner[19] */ 1'b0,
        /* cinner[18] */ |{ &{G[17]},
                            &{G[16], P[17]},
                            &{G[15], P[16], P[17]},
                            &{G[14], P[15], P[16], P[17]},
                            &{G[13], P[14], P[15], P[16], P[17]},
                            &{G[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], P[17], cin}},
        // /* cinner[18] */ 1'b0,
        /* cinner[17] */ |{ &{G[16]},
                            &{G[15], P[16]},
                            &{G[14], P[15], P[16]},
                            &{G[13], P[14], P[15], P[16]},
                            &{G[12], P[13], P[14], P[15], P[16]},
                            &{G[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], P[16], cin}},
        // /* cinner[17] */ 1'b0,
        /* cinner[16] */ |{ &{G[15]},
                            &{G[14], P[15]},
                            &{G[13], P[14], P[15]},
                            &{G[12], P[13], P[14], P[15]},
                            &{G[11], P[12], P[13], P[14], P[15]},
                            &{G[10], P[11], P[12], P[13], P[14], P[15]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14], P[15]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], P[15], cin}},
        // /* cinner[16] */ 1'b0,
        /* cinner[15] */ |{ &{G[14]},
                            &{G[13], P[14]},
                            &{G[12], P[13], P[14]},
                            &{G[11], P[12], P[13], P[14]},
                            &{G[10], P[11], P[12], P[13], P[14]},
                            &{G[ 9], P[10], P[11], P[12], P[13], P[14]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], P[14], cin}},
        // /* cinner[15] */ 1'b0,
        /* cinner[14] */ |{ &{G[13]},
                            &{G[12], P[13]},
                            &{G[11], P[12], P[13]},
                            &{G[10], P[11], P[12], P[13]},
                            &{G[ 9], P[10], P[11], P[12], P[13]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12], P[13]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], P[13], cin}},
        // /* cinner[14] */ 1'b0,
        /* cinner[13] */ |{ &{G[12]},
                            &{G[11], P[12]},
                            &{G[10], P[11], P[12]},
                            &{G[ 9], P[10], P[11], P[12]},
                            &{G[ 8], P[ 9], P[10], P[11], P[12]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11], P[12]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], P[12], cin}},
        // /* cinner[13] */ 1'b0,
        /* cinner[12] */ |{ &{G[11]},
                            &{G[10], P[11]},
                            &{G[ 9], P[10], P[11]},
                            &{G[ 8], P[ 9], P[10], P[11]},
                            &{G[ 7], P[ 8], P[ 9], P[10], P[11]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], P[11], cin}},
        // /* cinner[12] */ 1'b0,
        /* cinner[11] */ |{ &{G[10]},
                            &{G[ 9], P[10]},
                            &{G[ 8], P[ 9], P[10]},
                            &{G[ 7], P[ 8], P[ 9], P[10]},
                            &{G[ 6], P[ 7], P[ 8], P[ 9], P[10]},
                            &{G[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10]}, 
                            &{G[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10]}, 
                            &{G[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10]}, 
                            &{G[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10]},
                            &{G[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10]},
                            &{G[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10]},
                            &{P[ 0], P[ 1], P[ 2], P[ 3], P[ 4], P[ 5], P[ 6], P[ 7], P[ 8], P[ 9], P[10], cin}},
        // /* cinner[11] */ 1'b0,
        /* cinner[10] */ |{ &{G[9]},
                            &{G[8], P[9]},
                            &{G[7], P[8], P[9]},
                            &{G[6], P[7], P[8], P[9]},
                            &{G[5], P[6], P[7], P[8], P[9]}, 
                            &{G[4], P[5], P[6], P[7], P[8], P[9]}, 
                            &{G[3], P[4], P[5], P[6], P[7], P[8], P[9]}, 
                            &{G[2], P[3], P[4], P[5], P[6], P[7], P[8], P[9]},
                            &{G[1], P[2], P[3], P[4], P[5], P[6], P[7], P[8], P[9]},
                            &{G[0], P[1], P[2], P[3], P[4], P[5], P[6], P[7], P[8], P[9]},
                            &{P[0], P[1], P[2], P[3], P[4], P[5], P[6], P[7], P[8], P[9], cin}},
        // /* cinner[10] */ 1'b0,
        /* cinner[ 9] */ |{ &{G[8]},
                            &{G[7], P[8]},
                            &{G[6], P[7], P[8]},
                            &{G[5], P[6], P[7], P[8]}, 
                            &{G[4], P[5], P[6], P[7], P[8]}, 
                            &{G[3], P[4], P[5], P[6], P[7], P[8]}, 
                            &{G[2], P[3], P[4], P[5], P[6], P[7], P[8]},
                            &{G[1], P[2], P[3], P[4], P[5], P[6], P[7], P[8]},
                            &{G[0], P[1], P[2], P[3], P[4], P[5], P[6], P[7], P[8]},
                            &{P[0], P[1], P[2], P[3], P[4], P[5], P[6], P[7], P[8], cin}},
        // /* cinner[ 9] */ 1'b0,
        /* cinner[ 8] */ |{ &{G[7]},
                            &{G[6], P[7]},
                            &{G[5], P[6], P[7]}, 
                            &{G[4], P[5], P[6], P[7]}, 
                            &{G[3], P[4], P[5], P[6], P[7]}, 
                            &{G[2], P[3], P[4], P[5], P[6], P[7]},
                            &{G[1], P[2], P[3], P[4], P[5], P[6], P[7]},
                            &{G[0], P[1], P[2], P[3], P[4], P[5], P[6], P[7]},
                            &{P[0], P[1], P[2], P[3], P[4], P[5], P[6], P[7], cin}},
        // /* cinner[ 8] */ 1'b0,
        /* carry[ 7] */  |{ &{G[6]}, 
                            &{G[5], P[6]},
                            &{G[4], P[5], P[6]},
                            &{G[3], P[4], P[5], P[6]},
                            &{G[2], P[3], P[4], P[5], P[6]},
                            &{G[1], P[2], P[3], P[4], P[5], P[6]},
                            &{G[0], P[1], P[2], P[3], P[4], P[5], P[6]},
                            &{P[0], P[1], P[2], P[3], P[4], P[5], P[6], cin}},
        // /* cinner[ 7] */ 1'b0,
        /* cinner[ 6] */ |{ &{G[5]},
                            &{G[4], P[5]},
                            &{G[3], P[4], P[5]},
                            &{G[2], P[3], P[4], P[5]},
                            &{G[1], P[2], P[3], P[4], P[5]},
                            &{G[0], P[1], P[2], P[3], P[4], P[5]},
                            &{P[0], P[1], P[2], P[3], P[4], P[5] & cin}},
        // /* cinner[ 6] */ 1'b0
        /* cinner[ 5] */ |{ &{G[4]},
                            &{G[3], P[4]},
                            &{G[2], P[3], P[4]},
                            &{G[1], P[2], P[3], P[4]},
                            &{G[0], P[1], P[2], P[3], P[4]},
                            &{P[0], P[1], P[2], P[3], P[4] & cin}},
        // /* cinner[ 5] */ 1'b0,
        /* cinner[ 4] */ |{ &{G[3]},
                            &{G[2], P[3]},
                            &{G[1], P[2], P[3]},
                            &{G[0], P[1], P[2], P[3]},
                            &{P[0], P[1], P[2], P[3], cin}},
        // /* cinner[ 4] */ 1'b0,
        /* cinner[ 3] */ |{ &{G[2]},
                            &{G[1],P[2]},
                            &{G[0],P[1], P[2]},
                            &{P[0],P[1], P[2], cin}},
        // /* cinner[ 3] */ 1'b0,
        /* cinner[ 2] */ |{ &{G[1]},
                            &{G[0], P[1]},
                            &{P[0], P[1], cin}},
        // /* cinner[ 2] */ 1'b0, 
        /* cinner[ 1] */ |{ &{G[0]}, 
                            &{P[0],cin}},
        // /* cinner[ 1] */ 1'b0,
        /* cinner[ 0] */ |{ &{cin}}
        // /* cinner[ 0] */ 1'b0
    };

endmodule

module GrpPG(
    input  wire [31:0] op1,
    input  wire [31:0] op2,
    output wire [31:0] P,
    output wire [31:0] G
);

    ModP modP0( .op1(op1[0]), .op2(op2[0]), .P(P[0]) );
    ModG modG0( .op1(op1[0]), .op2(op2[0]), .G(G[0]) );

    ModP modP1( .op1(op1[1]), .op2(op2[1]), .P(P[1]) );
    ModG modG1( .op1(op1[1]), .op2(op2[1]), .G(G[1]) );

    ModP modP2( .op1(op1[2]), .op2(op2[2]), .P(P[2]) );
    ModG modG2( .op1(op1[2]), .op2(op2[2]), .G(G[2]) );

    ModP modP3( .op1(op1[3]), .op2(op2[3]), .P(P[3]) );
    ModG modG3( .op1(op1[3]), .op2(op2[3]), .G(G[3]) );

    ModP modP4( .op1(op1[4]), .op2(op2[4]), .P(P[4]) );
    ModG modG4( .op1(op1[4]), .op2(op2[4]), .G(G[4]) );

    ModP modP5( .op1(op1[5]), .op2(op2[5]), .P(P[5]) );
    ModG modG5( .op1(op1[5]), .op2(op2[5]), .G(G[5]) );

    ModP modP6( .op1(op1[6]), .op2(op2[6]), .P(P[6]) );
    ModG modG6( .op1(op1[6]), .op2(op2[6]), .G(G[6]) );

    ModP modP7( .op1(op1[7]), .op2(op2[7]), .P(P[7]) );
    ModG modG7( .op1(op1[7]), .op2(op2[7]), .G(G[7]) );

    ModP modP8( .op1(op1[8]), .op2(op2[8]), .P(P[8]) );
    ModG modG8( .op1(op1[8]), .op2(op2[8]), .G(G[8]) );

    ModP modP9( .op1(op1[9]), .op2(op2[9]), .P(P[9]) );
    ModG modG9( .op1(op1[9]), .op2(op2[9]), .G(G[9]) );

    ModP modP10( .op1(op1[10]), .op2(op2[10]), .P(P[10]) );
    ModG modG10( .op1(op1[10]), .op2(op2[10]), .G(G[10]) );

    ModP modP11( .op1(op1[11]), .op2(op2[11]), .P(P[11]) );
    ModG modG11( .op1(op1[11]), .op2(op2[11]), .G(G[11]) );

    ModP modP12( .op1(op1[12]), .op2(op2[12]), .P(P[12]) );
    ModG modG12( .op1(op1[12]), .op2(op2[12]), .G(G[12]) );

    ModP modP13( .op1(op1[13]), .op2(op2[13]), .P(P[13]) );
    ModG modG13( .op1(op1[13]), .op2(op2[13]), .G(G[13]) );

    ModP modP14( .op1(op1[14]), .op2(op2[14]), .P(P[14]) );
    ModG modG14( .op1(op1[14]), .op2(op2[14]), .G(G[14]) );

    ModP modP15( .op1(op1[15]), .op2(op2[15]), .P(P[15]) );
    ModG modG15( .op1(op1[15]), .op2(op2[15]), .G(G[15]) );

    ModP modP16( .op1(op1[16]), .op2(op2[16]), .P(P[16]) );
    ModG modG16( .op1(op1[16]), .op2(op2[16]), .G(G[16]) );

    ModP modP17( .op1(op1[17]), .op2(op2[17]), .P(P[17]) );
    ModG modG17( .op1(op1[17]), .op2(op2[17]), .G(G[17]) );

    ModP modP18( .op1(op1[18]), .op2(op2[18]), .P(P[18]) );
    ModG modG18( .op1(op1[18]), .op2(op2[18]), .G(G[18]) );

    ModP modP19( .op1(op1[19]), .op2(op2[19]), .P(P[19]) );
    ModG modG19( .op1(op1[19]), .op2(op2[19]), .G(G[19]) );

    ModP modP20( .op1(op1[20]), .op2(op2[20]), .P(P[20]) );
    ModG modG20( .op1(op1[20]), .op2(op2[20]), .G(G[20]) );

    ModP modP21( .op1(op1[21]), .op2(op2[21]), .P(P[21]) );
    ModG modG21( .op1(op1[21]), .op2(op2[21]), .G(G[21]) );

    ModP modP22( .op1(op1[22]), .op2(op2[22]), .P(P[22]) );
    ModG modG22( .op1(op1[22]), .op2(op2[22]), .G(G[22]) );

    ModP modP23( .op1(op1[23]), .op2(op2[23]), .P(P[23]) );
    ModG modG23( .op1(op1[23]), .op2(op2[23]), .G(G[23]) );

    ModP modP24( .op1(op1[24]), .op2(op2[24]), .P(P[24]) );
    ModG modG24( .op1(op1[24]), .op2(op2[24]), .G(G[24]) );

    ModP modP25( .op1(op1[25]), .op2(op2[25]), .P(P[25]) );
    ModG modG25( .op1(op1[25]), .op2(op2[25]), .G(G[25]) );

    ModP modP26( .op1(op1[26]), .op2(op2[26]), .P(P[26]) );
    ModG modG26( .op1(op1[26]), .op2(op2[26]), .G(G[26]) );

    ModP modP27( .op1(op1[27]), .op2(op2[27]), .P(P[27]) );
    ModG modG27( .op1(op1[27]), .op2(op2[27]), .G(G[27]) );

    ModP modP28( .op1(op1[28]), .op2(op2[28]), .P(P[28]) );
    ModG modG28( .op1(op1[28]), .op2(op2[28]), .G(G[28]) );

    ModP modP29( .op1(op1[29]), .op2(op2[29]), .P(P[29]) );
    ModG modG29( .op1(op1[29]), .op2(op2[29]), .G(G[29]) );

    ModP modP30( .op1(op1[30]), .op2(op2[30]), .P(P[30]) );
    ModG modG30( .op1(op1[30]), .op2(op2[30]), .G(G[30]) );

    ModP modP31( .op1(op1[31]), .op2(op2[31]), .P(P[31]) );
    ModG modG31( .op1(op1[31]), .op2(op2[31]), .G(G[31]) );

endmodule

module ModP(
    input  wire op1,
    input  wire op2,
    output wire P
);

    assign P = op1 ^ op2;

endmodule

module ModG(
    input  wire op1,
    input  wire op2,
    output wire G
);

    assign G = op1 & op2;

endmodule