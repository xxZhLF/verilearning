module Add64(
    input  wire [63:0] op1,
    input  wire [63:0] op2,
    output wire [63:0] sum
);



endmodule